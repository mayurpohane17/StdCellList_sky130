* SPICE3 file created from sky130_vsdinv_1x.ext - technology: sky130A

.option scale=0.01u

.subckt sky130_vsdinv_1x A Y VGND VPWR VPB
X0 Y A VGND VGND sky130_fd_pr__nfet_01v8 w=43 l=15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8 w=70 l=15
C0 Y VPB 0.00fF
C1 VPWR A 0.01fF
C2 Y A 0.03fF
C3 VPWR VPB 0.02fF
C4 Y VPWR 0.07fF
C5 Y VGND 0.18fF
C6 VPWR VGND 0.23fF
C7 VPB VGND 0.15fF
.ends
